--===========================================================
--     ___        _      __   ____                         
--    /   |_   __(____  / /  / __ )_________ _      ______ 
--   / /| | | / / / _ \/ /  / __  / ___/ __ | | /| / / __ \
--  / ___ | |/ / /  __/ /  / /_/ / /  / /_/ | |/ |/ / / / /
-- /_/  |_|___/_/\___/_/  /_____/_/   \____/|__/|__/_/ /_/ 
--===========================================================
-- Advanced Logic Design	
-- Assignment 1
--===========================================================

entity demux is

	port(
	
		x, B, A : in bit;
		D0, D1, D2, D3 : out bit
		
);

end entity;



architecture demux_arc of demux is
begin

	D0 <= (x) and ((not B) and (not A));
	D1 <= (x) and ((not B) and (A));
	D2 <= (x) and ((B) and (not A));
	D3 <= (x) and ((B) and (A));
	
end demux_arc;
